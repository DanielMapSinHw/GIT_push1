version https://git-lfs.github.com/spec/v1
oid sha256:d42bade6c7a1c57910c1a852482e003110151615682c5457eafc3d7b71ff2f38
size 836
